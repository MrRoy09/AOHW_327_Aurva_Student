`timescale 1ns / 1ps

`define N 256
`define Q 132120577
`define K 27
`define barret_const 136348167

